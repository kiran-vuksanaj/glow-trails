`timescale 1ns / 1ps
`default_nettype none

module memory
  #(
    parameter WIDTH = 240)
   (
    input wire row,
    input wire column,
    output logic valid,
	output logic app_addr_mt
	);
   // your code here
	
	
	
	
endmodule


`default_nettype wire

